module lab_002_partb (
  input A,
  input B,
  input C,
  output F
);

  /* put your variable declarations here */


  /* put your gate instances here */

endmodule
