module lab_003_parta (
  input A, B, C,
  output G
);

endmodule
