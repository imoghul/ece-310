module lab_003_partc (
  input A, B, C, D,
  output F
);

endmodule
